//=========================================================================
// 5-Stage Simple Pipelined Processor
//=========================================================================

`ifndef LAB2_PROC_PIPELINED_PROC_BASE_V
`define LAB2_PROC_PIPELINED_PROC_BASE_V

`include "vc/mem-msgs.v"
`include "vc/queues.v"
`include "vc/trace.v"

`include "lab2_proc/TinyRV2InstVRTL.v"
`include "lab2_proc/ProcBaseCtrlVRTL.v"
`include "lab2_proc/ProcBaseDpathVRTL.v"
`include "lab2_proc/DropUnitVRTL.v"

module lab2_proc_ProcBaseVRTL
#(
  parameter p_num_cores = 1
)
(
  input  logic         clk,
  input  logic         reset,

  // core_id is an input port rather than a parameter so that
  // the module only needs to be compiled once. If it were a parameter,
  // each core would be compiled separately.
  input  logic [31:0]  core_id,

  // From mngr streaming port

  input  logic [31:0]  mngr2proc_msg,
  input  logic         mngr2proc_val,
  output logic         mngr2proc_rdy,

  // To mngr streaming port

  output logic [31:0]  proc2mngr_msg,
  output logic         proc2mngr_val,
  input  logic         proc2mngr_rdy,

  // Instruction Memory Request Port

  output mem_req_4B_t  imemreq_msg,
  output logic         imemreq_val,
  input  logic         imemreq_rdy,

  // Instruction Memory Response Port

  input  mem_resp_4B_t imemresp_msg,
  input  logic         imemresp_val,
  output logic         imemresp_rdy,

  // Data Memory Request Port

  output mem_req_4B_t  dmemreq_msg,
  output logic         dmemreq_val,
  input  logic         dmemreq_rdy,

  // Data Memory Response Port

  input  mem_resp_4B_t dmemresp_msg,
  input  logic         dmemresp_val,
  output logic         dmemresp_rdy,

  // stats output

  output logic         commit_inst,

  output logic         stats_en
 // output logic         inst_X_direct

);

  //----------------------------------------------------------------------
  // data mem req/resp
  //----------------------------------------------------------------------

  // imemreq before pack

  logic [31:0] imemreq_msg_addr;

  // imemreq_enq signals after pack before bypass queue

  mem_req_4B_t imemreq_enq_msg;
  logic        imemreq_enq_val;
  logic        imemreq_enq_rdy;

  // dmem req before pack

  logic [31:0] dmemreq_msg_addr;

  // dmemreq after pack before bypass queue

  mem_req_4B_t dmemreq_enq_msg;
  logic        dmemreq_enq_val;
  logic        dmemreq_enq_rdy;
  logic [31:0] dmemreq_msg_data;

  // proc2mngr signals before bypass queue

  logic [31:0] proc2mngr_enq_msg;
  logic        proc2mngr_enq_val;
  logic        proc2mngr_enq_rdy;

  // imemresp signals after the drop unit

  logic        imemresp_val_drop;
  logic        imemresp_rdy_drop;

  // imemresp drop signal

  logic        imemresp_drop;

  // control signals (ctrl->dpath)

  logic        reg_en_F;
  logic [1:0]  pc_sel_F;

  logic        reg_en_D;
  logic        op1_sel_D;
  logic [1:0]  op2_sel_D;
  logic [1:0]  csrr_sel_D;
  logic [2:0]  imm_type_D;

  logic        reg_en_X;
  logic [3:0]  alu_fn_X;
  logic [1:0]  ex_result_sel_X;

  logic        reg_en_M;
  logic        wb_result_sel_M;

  logic        reg_en_W;
  logic [4:0]  rf_waddr_W;
  logic        rf_wen_W;
  logic        stats_en_wen_W;

  // status signals (dpath->ctrl)

  logic [31:0] inst_D;
  logic        br_cond_eq_X;
  logic        br_cond_lt_X;
  logic        br_cond_ltu_X;
  
  //here
  logic [31:0] rf_rdata0_D;
  logic [31:0] rf_rdata1_D;
  logic [31:0] alu_result_X;
  logic [31:0] op1_X;
  logic [31:0] op2_X;  
  logic [31:0] ex_result_M;
  logic [31:0] wb_result_W; 
  logic [31:0] ex_result_X;
  logic [31:0] imm_D;
  logic [31:0] jal_target_D;
  logic [31:0] imul_resp_msg;
  
  /// testing only
  logic         inst_X_direct;
  logic         osquash_D;
  //----------------------------------------------------------------------
  // Pack Memory Request Messages
  //----------------------------------------------------------------------
  
  assign imemreq_enq_msg.type_  = `VC_MEM_REQ_MSG_TYPE_READ;
  assign imemreq_enq_msg.opaque = 8'b0;
  assign imemreq_enq_msg.addr   = imemreq_msg_addr;
  assign imemreq_enq_msg.len    = 2'd0;
  assign imemreq_enq_msg.data   = 32'bx;
  
  always_comb begin
    if (inst_X_direct==1) begin
         dmemreq_enq_msg.type_  = `VC_MEM_REQ_MSG_TYPE_WRITE;   
         dmemreq_enq_msg.opaque = 8'b0;
         dmemreq_enq_msg.addr   = dmemreq_msg_addr;
         dmemreq_enq_msg.len    = 2'd0;
         dmemreq_enq_msg.data   = dmemreq_msg_data;
    end
    else begin
         dmemreq_enq_msg.type_  = `VC_MEM_REQ_MSG_TYPE_READ;
         dmemreq_enq_msg.opaque = 8'b0;
         dmemreq_enq_msg.addr   = dmemreq_msg_addr;
         dmemreq_enq_msg.len    = 2'd0;
         dmemreq_enq_msg.data   = 32'b0;
    end
  end

  //----------------------------------------------------------------------
  // Imem Drop Unit
  //----------------------------------------------------------------------

  mem_resp_4B_t imemresp_msg_drop;

  vc_DropUnit #($bits(mem_resp_4B_t)) imem_drop_unit
  (
    .clk      (clk),
    .reset    (reset),

    .drop     (imemresp_drop),

    .in_msg   (imemresp_msg),
    .in_val   (imemresp_val),
    .in_rdy   (imemresp_rdy),

    .out_msg  (imemresp_msg_drop),
    .out_val  (imemresp_val_drop),
    .out_rdy  (imemresp_rdy_drop)
  );

  //----------------------------------------------------------------------
  // Control UnitRS2
  //----------------------------------------------------------------------
  logic        imul_req_rdy_D;
  logic        imul_req_val_D;
  logic        imul_resp_val_X;
  logic        imul_resp_rdy_X;
  
  lab2_proc_ProcBaseCtrlVRTL ctrl
  (
    .clk                    (clk),
    .reset                  (reset),

    // Instruction Memory Port

    .imemreq_val            (imemreq_enq_val),
    .imemreq_rdy            (imemreq_enq_rdy),
    .imemresp_val           (imemresp_val_drop),
    .imemresp_rdy           (imemresp_rdy_drop),
    .imul_req_val_D         (imul_req_val_D),// we add this input of imul
    .imul_resp_val_X        (imul_resp_val_X),// we add this input of imul
    .imul_req_rdy_D         (imul_req_rdy_D),//we add this output of l
    .imul_resp_rdy_X        (imul_resp_rdy_X),

    // Drop signal

    .imemresp_drop          (imemresp_drop),

    // Data Memory Port

    .dmemreq_val            (dmemreq_enq_val),
    .dmemreq_rdy            (dmemreq_enq_rdy),
    .dmemresp_val           (dmemresp_val),
    .dmemresp_rdy           (dmemresp_rdy),

    // mngr communication ports

    .mngr2proc_val          (mngr2proc_val),
    .mngr2proc_rdy          (mngr2proc_rdy),
    .proc2mngr_val          (proc2mngr_enq_val),
    .proc2mngr_rdy          (proc2mngr_enq_rdy),

    // control signals (ctrl->dpath)

    .reg_en_F               (reg_en_F),
    .pc_sel_F               (pc_sel_F),

    .reg_en_D               (reg_en_D),
    .op1_sel_D              (op1_sel_D),
    .op2_sel_D              (op2_sel_D),
    .csrr_sel_D             (csrr_sel_D),
    .imm_type_D             (imm_type_D),

    .reg_en_X               (reg_en_X),
    .alu_fn_X               (alu_fn_X),

    .reg_en_M               (reg_en_M),
    .wb_result_sel_M        (wb_result_sel_M),

    .reg_en_W               (reg_en_W),
    .rf_waddr_W             (rf_waddr_W),
    .rf_wen_W               (rf_wen_W),
    .stats_en_wen_W         (stats_en_wen_W),

    // status signals (dpath->ctrl)

    .inst_D                 (inst_D),
    .br_cond_eq_X           (br_cond_eq_X),
    .br_cond_lt_X           (br_cond_lt_X),
    .br_cond_ltu_X          (br_cond_ltu_X),
    .ex_result_sel_X        (ex_result_sel_X),

    .commit_inst            (commit_inst),
    .inst_X_direct          (inst_X_direct),
    .osquash_D              (osquash_D)             
  );

  //----------------------------------------------------------------------
  // Bypass Queue
  //----------------------------------------------------------------------

  logic [1:0] imem_queue_num_free_entries;

  vc_Queue#(`VC_QUEUE_BYPASS,$bits(mem_req_4B_t),2) imem_queue
  (
    .clk     (clk),
    .reset   (reset),
    .num_free_entries(imem_queue_num_free_entries),
    .enq_val (imemreq_enq_val),
    .enq_rdy (imemreq_enq_rdy),
    .enq_msg (imemreq_enq_msg),
    .deq_val (imemreq_val),
    .deq_rdy (imemreq_rdy),
    .deq_msg (imemreq_msg)
  );

  logic dmem_queue_num_free_entries;

  vc_Queue#(`VC_QUEUE_BYPASS,$bits(mem_req_4B_t),1) dmem_queue
  (
    .clk     (clk),
    .reset   (reset),
    .num_free_entries(dmem_queue_num_free_entries),
    .enq_val (dmemreq_enq_val),
    .enq_rdy (dmemreq_enq_rdy),
    .enq_msg (dmemreq_enq_msg),
    .deq_val (dmemreq_val),
    .deq_rdy (dmemreq_rdy),
    .deq_msg (dmemreq_msg)
  );

  logic proc2mngr_queue_num_free_entries;

  vc_Queue#(`VC_QUEUE_BYPASS,32,1) proc2mngr_queue
  (
    .clk     (clk),
    .reset   (reset),
    .num_free_entries(proc2mngr_queue_num_free_entries),
    .enq_val (proc2mngr_enq_val),
    .enq_rdy (proc2mngr_enq_rdy),
    .enq_msg (proc2mngr_enq_msg),
    .deq_val (proc2mngr_val),
    .deq_rdy (proc2mngr_rdy),
    .deq_msg (proc2mngr_msg)
  );

  //----------------------------------------------------------------------
  // Datapath
  //----------------------------------------------------------------------
  
  lab2_proc_ProcBaseDpathVRTL
  #(
    .p_num_cores             (p_num_cores)
  )
  dpath
  (
    .clk                     (clk),
    .reset                   (reset),
    .imul_req_val_D          (imul_req_val_D),// we add this input of imul
    .imul_resp_val_X         (imul_resp_val_X),// we add this input of imul
    .imul_req_rdy_D          (imul_req_rdy_D),//we add this output of l
    .imul_resp_rdy_X         (imul_resp_rdy_X),//we add this output of imul  

    // core id
    .core_id                 (core_id),

    // Instruction Memory Port

    .imemreq_msg_addr        (imemreq_msg_addr),
    .imemresp_msg            (imemresp_msg_drop),
    //.dmemreq_msg_data        (dmemreq_msg_data),
    // Data Memory Port

    .dmemreq_msg_addr        (dmemreq_msg_addr),
    .dmemresp_msg_data       (dmemresp_msg.data),
    .dmemreq_msg_data        (dmemreq_msg_data),
    // mngr communication ports

    .mngr2proc_data          (mngr2proc_msg),
    .proc2mngr_data          (proc2mngr_enq_msg),

    // control signals (ctrl->dpath)

    .imemresp_val_drop       (imemresp_val_drop),
    .imemresp_rdy_drop       (imemresp_rdy_drop),
    .imemresp_drop           (imemresp_drop),

    .reg_en_F                (reg_en_F),
    .pc_sel_F                (pc_sel_F),

    .reg_en_D                (reg_en_D),
    .op1_sel_D               (op1_sel_D),
    .op2_sel_D               (op2_sel_D),
    .csrr_sel_D              (csrr_sel_D),
    .imm_type_D              (imm_type_D),

    .reg_en_X                (reg_en_X),
    .alu_fn_X                (alu_fn_X),

    .reg_en_M                (reg_en_M),
    .wb_result_sel_M         (wb_result_sel_M),

    .reg_en_W                (reg_en_W),
    .rf_waddr_W              (rf_waddr_W),
    .rf_wen_W                (rf_wen_W),
    .stats_en_wen_W          (stats_en_wen_W),
    .ex_result_sel_X         (ex_result_sel_X),
    .imul_resp_msg           (imul_resp_msg),
    // status signals (dpath->ctrl)

    .inst_D                  (inst_D),
    .br_cond_eq_X            (br_cond_eq_X),
    .br_cond_lt_X           (br_cond_lt_X),
    .br_cond_ltu_X          (br_cond_ltu_X),

    // stats_en

    .stats_en                (stats_en),
    .rf_rdata0_D             (rf_rdata0_D),
    .rf_rdata1_D             (rf_rdata1_D),
    .alu_result_X            (alu_result_X),
    .op1_X                   (op1_X),
    .op2_X                   (op2_X),
    .ex_result_M             (ex_result_M),
    .wb_result_W             (wb_result_W),
    .ex_result_X             (ex_result_X),
    .imm_D                   (imm_D),
    .jal_target_D            (jal_target_D)
  );

  //----------------------------------------------------------------------
  // Line tracing
  //----------------------------------------------------------------------

  `ifndef SYNTHESIS

  rv2isa_InstTasks rv2isa();

  logic [`VC_TRACE_NBITS-1:0] str;
  `VC_TRACE_BEGIN
  begin

    if ( !ctrl.val_F )
      vc_trace.append_chars( trace_str, " ", 8 );
    else if ( ctrl.squash_F ) begin
      vc_trace.append_str( trace_str, "~" );
      vc_trace.append_chars( trace_str, " ", 8-1 );
    end else if ( ctrl.stall_F ) begin
      vc_trace.append_str( trace_str, "#" );
      vc_trace.append_chars( trace_str, " ", 8-1 );
    end else begin
      $sformat( str, "%x", dpath.pc_F );
      vc_trace.append_str( trace_str, str );
    end

    vc_trace.append_str( trace_str, "|" );

    if ( !ctrl.val_D )
      vc_trace.append_chars( trace_str, " ", 23 );
    else if ( ctrl.squash_D ) begin
      vc_trace.append_str( trace_str, "~" );
      vc_trace.append_chars( trace_str, " ", 23-1 );
    end else if ( ctrl.stall_D ) begin
      vc_trace.append_str( trace_str, "#" );
      vc_trace.append_chars( trace_str, " ", 23-1 );
    end else
      vc_trace.append_str( trace_str, { 3896'b0, rv2isa.disasm( ctrl.inst_D ) } );

    vc_trace.append_str( trace_str, "|" );

    if ( !ctrl.val_X )
      vc_trace.append_chars( trace_str, " ", 4 );
    else if ( ctrl.stall_X ) begin
      vc_trace.append_str( trace_str, "#" );
      vc_trace.append_chars( trace_str, " ", 4-1 );
    end else
      vc_trace.append_str( trace_str, { 4064'b0, rv2isa.disasm_tiny( ctrl.inst_X ) } );
     
    if ( !ctrl.val_M )
      vc_trace.append_chars( trace_str, " ", 4 );
    else if ( ctrl.stall_M ) begin
      vc_trace.append_str( trace_str, "#" );
      vc_trace.append_chars( trace_str, " ", 4-1 );
    end else
      vc_trace.append_str( trace_str, { 4064'b0, rv2isa.disasm_tiny( ctrl.inst_M ) } );

    vc_trace.append_str( trace_str, "|" );

    if ( !ctrl.val_W )
      vc_trace.append_chars( trace_str, " ", 4 );
    else if ( ctrl.stall_W ) begin
      vc_trace.append_str( trace_str, "#" );
      vc_trace.append_chars( trace_str, " ", 4-1 );
    end else
      vc_trace.append_str( trace_str, { 4064'b0, rv2isa.disasm_tiny( ctrl.inst_W ) } );
    //testing only  
    //vc_trace.append_str( trace_str, "| machine code:" );  
    // $sformat( str, "%x", dpath.inst_D  );
   // vc_trace.append_str( trace_str, str );
   vc_trace.append_str( trace_str, "| pc_sel:" );  
     $sformat( str, "%x",pc_sel_F);
    vc_trace.append_str( trace_str, str );
    /*
    vc_trace.append_str( trace_str, "| osquash:" );  
     $sformat( str, "%x", osquash_D);
    vc_trace.append_str( trace_str, str );
    */
   vc_trace.append_str( trace_str, "| imm:" );  
     $sformat( str, "%x", dpath.imm_D);
    vc_trace.append_str( trace_str, str );
   /* 
    vc_trace.append_str( trace_str, "| jal_target_D ");  
     $sformat( str, "%x", dpath.jal_target_D);
    vc_trace.append_str( trace_str, str );
    */
    /*    
    vc_trace.append_str( trace_str, "| RS1:" );  
     $sformat( str, "%x", dpath.rf_rdata0_D );
    vc_trace.append_str( trace_str, str );
    
     vc_trace.append_str( trace_str, "| RS2:" );  
     $sformat( str, "%x", dpath.rf_rdata1_D );
    vc_trace.append_str( trace_str, str );
    */
    vc_trace.append_str( trace_str, "| RS2:" );  
     $sformat( str, "%x", dpath.rf_rdata1_D );
    vc_trace.append_str( trace_str, str );
    /*
    vc_trace.append_str( trace_str, "| val_D:" );  
     $sformat( str, "%x", imul_req_val_D);
    vc_trace.append_str( trace_str, str );
    
    vc_trace.append_str( trace_str, "| rdy_D:" );  
     $sformat( str, "%x", imul_req_rdy_D);
    vc_trace.append_str( trace_str, str );
    
    vc_trace.append_str( trace_str, "| val_X:" );  
     $sformat( str, "%x", imul_resp_val_X);
    vc_trace.append_str( trace_str, str );
    
    vc_trace.append_str( trace_str, "| rdy_X:" );  
     $sformat( str, "%x", imul_resp_rdy_X);
    vc_trace.append_str( trace_str, str );
    
    vc_trace.append_str( trace_str, "| OP2:" );  
     $sformat( str, "%x", dpath.op2_X);
    vc_trace.append_str( trace_str, str );
    */
     vc_trace.append_str( trace_str, "| ALU_Out:" );  
     $sformat( str, "%x", dpath.alu_result_X);
    vc_trace.append_str( trace_str, str );
    /*
    vc_trace.append_str( trace_str, "| msg:" );  
     $sformat( str, "%x", dpath.imul_resp_msg);
    vc_trace.append_str( trace_str, str );
    
    vc_trace.append_str( trace_str, "| br_cond_lt_X:" );  
     $sformat( str, "%x", br_cond_lt_X);
    vc_trace.append_str( trace_str, str );
    */
    /*
    vc_trace.append_str( trace_str, "| br_cond_eq:" );  
     $sformat( str, "%x", br_cond_eq_X);
    vc_trace.append_str( trace_str, str );
    */
    /*
    vc_trace.append_str( trace_str, "| dmemreq:" );  
     $sformat( str, "%x", dmemreq_msg_data);
    vc_trace.append_str( trace_str, str );
    
     vc_trace.append_str( trace_str, "| SW?=:" );  
     $sformat( str, "%x", inst_X_direct);
    vc_trace.append_str( trace_str, str );
    */
    /*
     vc_trace.append_str( trace_str, "| ex_result_sel_X:" );  
     $sformat( str, "%x", dpath. ex_result_sel_X);
    vc_trace.append_str( trace_str, str );
    
    vc_trace.append_str( trace_str, "ex_result_x:" );  
     $sformat( str, "%x", dpath.ex_result_X);
    vc_trace.append_str( trace_str, str );
    
    vc_trace.append_str( trace_str, "| wb_result_sel_M:" );  
     $sformat( str, "%x", dpath.wb_result_sel_M);
    vc_trace.append_str( trace_str, str );
    
    vc_trace.append_str( trace_str, "| ex_result_M:" );  
     $sformat( str, "%x", dpath.ex_result_M);
    vc_trace.append_str( trace_str, str );
    
    
    vc_trace.append_str( trace_str, "| Wb_result_W:" );  
     $sformat( str, "%x", dpath.wb_result_W);
    vc_trace.append_str( trace_str, str );
    
      vc_trace.append_str( trace_str, "| rf_wen_W:" );  
     $sformat( str, "%x", dpath.rf_wen_W);
    vc_trace.append_str( trace_str, str );
    */
     
  end
  `VC_TRACE_END

  vc_MemReqMsg4BTrace imemreq_trace
  (
    .clk   (clk),
    .reset (reset),
    .val   (imemreq_val),
    .rdy   (imemreq_rdy),
    .msg   (imemreq_msg)
  );

  vc_MemReqMsg4BTrace dmemreq_trace
  (
    .clk   (clk),
    .reset (reset),
    .val   (dmemreq_val),
    .rdy   (dmemreq_rdy),
    .msg   (dmemreq_msg)
  );

  vc_MemRespMsg4BTrace imemresp_trace
  (
    .clk   (clk),
    .reset (reset),
    .val   (imemresp_val),
    .rdy   (imemresp_rdy),
    .msg   (imemresp_msg)
  );

  vc_MemRespMsg4BTrace dmemresp_trace
  (
    .clk   (clk),
    .reset (reset),
    .val   (dmemresp_val),
    .rdy   (dmemresp_rdy),
    .msg   (dmemresp_msg)
  );

  `endif

endmodule

`endif

